----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:33:04 10/16/2018 
-- Design Name: 
-- Module Name:    FrBuf - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity FrBuf is
    Port ( next_col : in  STD_LOGIC_VECTOR (9 downto 0);
           row : in  STD_LOGIC_VECTOR (9 downto 0);
           pixel : out  STD_LOGIC;
           clk : in  STD_LOGIC);
end FrBuf;

architecture Behavioral of FrBuf is

signal mem_out, pixel_vec : unsigned(19 downto 0);
signal word_col : unsigned(4 downto 0);
signal address : unsigned(13 downto 0);
signal load : boolean; 
signal ncol, nrow: integer;


type framebuf_type is array (0 to 16383) of std_logic_vector(19 downto 0);
constant framebuffer: framebuf_type := (
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 0
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 1
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 2
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 3
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 4
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 5
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 6
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 7
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 8
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 9
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 10
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 11
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 12
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 13
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 14
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 15
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 16
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 17
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 18
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 19
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 20
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 21
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 22
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 23
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 24
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 25
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 26
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 27
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 28
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 29
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 30
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 31
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 32
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 33
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 34
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 35
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 36
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 37
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 38
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 39
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 40
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 41
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 42
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 43
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 44
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 45
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 46
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 47
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 48
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 49
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 50
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 51
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 52
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 53
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 54
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 55
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 56
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 57
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 58
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 59
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 60
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 61
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 62
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 63
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 64
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 65
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 66
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 67
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 68
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 69
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 70
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 71
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 72
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 73
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 74
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 75
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 76
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 77
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 78
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 79
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 80
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 81
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 82
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 83
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 84
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 85
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 86
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 87
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 88
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 89
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 90
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 91
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 92
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 93
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 94
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 95
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 96
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 97
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 98
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 99
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 100
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 101
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 102
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 103
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 104
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 105
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 106
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 107
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 108
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 109
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 110
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 111
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 112
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 113
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 114
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 115
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 116
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 117
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 118
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 119
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 120
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 121
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 122
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 123
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 124
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 125
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 126
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 127
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 128
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 129
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 130
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 131
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 132
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 133
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 134
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 135
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 136
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 137
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 138
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 139
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 140
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 141
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 142
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 143
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 144
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 145
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 146
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 147
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 148
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 149
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 150
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 151
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 152
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 153
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 154
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 155
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 156
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 157
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 158
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 159
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 160
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 161
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 162
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 163
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 164
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 165
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 166
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 167
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 168
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 169
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 170
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 171
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 172
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 173
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 174
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 175
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 176
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 177
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 178
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 179
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 180
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 181
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 182
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 183
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 184
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 185
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 186
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 187
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 188
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 189
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 190
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 191
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 192
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 193
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 194
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 195
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 196
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 197
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 198
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 199
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 200
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 201
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 202
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 203
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 204
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 205
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 206
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 207
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 208
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 209
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 210
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 211
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 212
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 213
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 214
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 215
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 216
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 217
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 218
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 219
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 220
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 221
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 222
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 223
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 224
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 225
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 226
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 227
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 228
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 229
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 230
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 231
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 232
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 233
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 234
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 235
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 236
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 237
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 238
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 239
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 240
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 241
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 242
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 243
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 244
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 245
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 246
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 247
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 248
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 249
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 250
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 251
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 252
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 253
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 254
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 255
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 256
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 257
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 258
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 259
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 260
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 261
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 262
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 263
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 264
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 265
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 266
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 267
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 268
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 269
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 270
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 271
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 272
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 273
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 274
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 275
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 276
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 277
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 278
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 279
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 280
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 281
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 282
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 283
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 284
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 285
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 286
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 287
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 288
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 289
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 290
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 291
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 292
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 293
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 294
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 295
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 296
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 297
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 298
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 299
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 300
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 301
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 302
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 303
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 304
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 305
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 306
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 307
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 308
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 309
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 310
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 311
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 312
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 313
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 314
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 315
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 316
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 317
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 318
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 319
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 320
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 321
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 322
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 323
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 324
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 325
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 326
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 327
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 328
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 329
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 330
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 331
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 332
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 333
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 334
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 335
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 336
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 337
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 338
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 339
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 340
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 341
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 342
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 343
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 344
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 345
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 346
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 347
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"02000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 348
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"06000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 349
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"07000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 350
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"07000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 351
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"0F000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 352
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"0F000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 353
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"0F800",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 354
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"0F800",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 355
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"1F800",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 356
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"7FF00",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 357
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"7FF00",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 358
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"FFF00",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 359
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFF80",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 360
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 361
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 362
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 363
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 364
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 365
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 366
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 367
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 368
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 369
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 370
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 371
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 372
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 373
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 374
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"10000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 375
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"10000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 376
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"10000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 377
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"10000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 378
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"10000",X"00000",X"00000",X"00003",X"FFFE0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 379
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"10000",X"00000",X"00000",X"00003",X"FFFF0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 380
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"10000",X"00000",X"00000",X"00003",X"FFFF0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 381
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"10000",X"00000",X"00000",X"00003",X"FFFF0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 382
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00003",X"FFFF0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 383
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00003",X"FFFF0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 384
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00003",X"FFFF0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 385
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 386
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 387
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 388
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 389
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"1FFFE",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 390
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 391
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 392
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 393
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 394
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 395
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"18000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 396
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"3C000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"00000",X"00400",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 397
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"3C000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"00000",X"00400",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 398
X"00000",X"00200",X"00000",X"00000",X"00000",X"00000",X"FF000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"00000",X"00400",X"00000",
X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 399
X"00000",X"00700",X"00000",X"00000",X"00000",X"00001",X"FF000",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"00000",X"00400",X"00000",
X"00200",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 400
X"00000",X"00600",X"00000",X"00000",X"00000",X"00001",X"FF800",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"00000",X"00400",X"00000",
X"00200",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 401
X"00000",X"00E00",X"00000",X"00000",X"00000",X"00001",X"FF800",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"00000",X"00400",X"00000",
X"00300",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 402
X"00000",X"00F80",X"00000",X"00000",X"00000",X"00001",X"FF800",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"3FFFF",X"FEE00",X"00000",
X"00300",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 403
X"00000",X"00F80",X"00000",X"00000",X"00000",X"00001",X"FF800",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"3FFFF",X"FFE00",X"00000",
X"00700",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 404
X"00000",X"00F00",X"00000",X"00000",X"00000",X"00001",X"FF800",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"3FFFF",X"FFF00",X"00000",
X"00780",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 405
X"00000",X"00600",X"00000",X"00000",X"00000",X"00003",X"FFC00",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"3FFFF",X"FFF00",X"00000",
X"00780",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 406
X"00000",X"00600",X"00000",X"00000",X"00000",X"00003",X"FFC00",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"3FFFF",X"FFF00",X"00000",
X"00FE0",X"00000",X"00000",X"00000",X"007FE",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 407
X"00000",X"00700",X"00000",X"00000",X"00000",X"00003",X"FFC00",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"3FFFF",X"FFF80",X"00000",
X"00FE0",X"00000",X"00000",X"00001",X"FCFFF",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 408
X"00000",X"00700",X"00000",X"00000",X"00000",X"00003",X"FFC00",X"00000",X"00000",X"00007",X"FFFF0",
X"00000",X"00000",X"00000",X"3FFFF",X"00000",X"00000",X"00000",X"00000",X"3FFFF",X"FFFC0",X"00000",
X"3FFF0",X"00000",X"00000",X"00001",X"FFFFF",X"00000",X"00000",X"00000",X"00000",X"00000",-- row 409
X"00000",X"00700",X"00000",X"00000",X"00000",X"00003",X"FFC00",X"00000",X"00000",X"00007",X"FFFF8",
X"00000",X"00000",X"00000",X"3FFFF",X"001FF",X"FFF00",X"00000",X"00000",X"3FFFF",X"FFFC0",X"00000",
X"3FFF0",X"00000",X"00000",X"0003F",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 410
X"00000",X"00300",X"00000",X"00000",X"00000",X"00003",X"FFC00",X"00000",X"00000",X"00007",X"FFFF8",
X"00000",X"00000",X"00000",X"3FFFF",X"00FFF",X"FFF00",X"00000",X"00000",X"3FFFF",X"FFFC0",X"00000",
X"7FFF0",X"00000",X"00000",X"000FF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 411
X"00000",X"00300",X"00000",X"00000",X"00000",X"00003",X"FFC00",X"00000",X"00000",X"00007",X"FFFF8",
X"00000",X"00000",X"00000",X"3FFFF",X"00FFF",X"FFF00",X"00000",X"00000",X"3FFFF",X"FFFC0",X"00000",
X"FFFF0",X"00000",X"00000",X"000FF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 412
X"00000",X"00300",X"00000",X"00000",X"00000",X"00003",X"FFC00",X"00000",X"00000",X"00007",X"FFFF8",
X"00000",X"00000",X"00000",X"7FFFF",X"00FFF",X"FFF00",X"00000",X"00000",X"3FFFF",X"FFFC0",X"00001",
X"FFFF0",X"00000",X"00000",X"000FF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 413
X"00000",X"00382",X"00000",X"00000",X"00000",X"00003",X"FFC00",X"00000",X"3C000",X"00007",X"FFFF8",
X"00000",X"00000",X"0003F",X"FFFFF",X"00FFF",X"FFF00",X"00000",X"00000",X"3FFFF",X"FFFC0",X"00003",
X"FFFF0",X"00000",X"00000",X"000FF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 414
X"00000",X"00392",X"20000",X"00000",X"00000",X"00003",X"FFC03",X"FFF80",X"7E000",X"00007",X"FFFFF",
X"FF000",X"00000",X"0003F",X"FFFFF",X"00FFF",X"FFF00",X"00000",X"01F80",X"3FFFF",X"FFFE0",X"0000F",
X"FFFF0",X"00000",X"00000",X"000FF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 415
X"00000",X"003CA",X"48000",X"00000",X"00000",X"00003",X"FFC07",X"FFF80",X"FF800",X"00007",X"FFFFF",
X"FF000",X"00000",X"0003F",X"FFFFF",X"00FFF",X"FFF00",X"00000",X"01F80",X"3FFFF",X"FFFE0",X"00007",
X"FFFF0",X"00000",X"00000",X"000FF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 416
X"00000",X"00387",X"80000",X"00000",X"00000",X"00003",X"FFC07",X"FFF83",X"FFE00",X"00007",X"FFFFF",
X"FF000",X"00000",X"0003F",X"FFFFF",X"00FFF",X"FFF00",X"00000",X"01F80",X"3FFFF",X"FFFE0",X"00007",
X"FFFF0",X"00000",X"00000",X"000FF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 417
X"00000",X"001FF",X"F0000",X"00000",X"00000",X"00003",X"FFC07",X"FFF87",X"FFE00",X"00007",X"FFFFF",
X"FF000",X"00000",X"0003F",X"FFFFF",X"00FFF",X"FFF00",X"00000",X"01F80",X"3FFFF",X"FFFE0",X"00007",
X"FFFF0",X"00000",X"00000",X"000FF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 418
X"00000",X"001CF",X"C0000",X"00000",X"00000",X"00003",X"FFC07",X"FFF87",X"FFF00",X"00007",X"FFFFF",
X"FF000",X"00000",X"0003F",X"FFFFF",X"00FFF",X"FFF00",X"00000",X"01F80",X"3FFFF",X"FFFE0",X"00007",
X"FFFF0",X"00F80",X"00000",X"000FF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 419
X"00000",X"001EF",X"C0000",X"00000",X"00000",X"00003",X"FFC07",X"FFF8F",X"FFF0F",X"80007",X"FFFFF",
X"FF000",X"00000",X"0003F",X"FFFFF",X"00FFF",X"FFF00",X"00000",X"01F80",X"3FFFF",X"FFFE0",X"00007",
X"FFFF0",X"01FE0",X"00000",X"000FF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 420
X"00000",X"001EF",X"C0000",X"00000",X"00000",X"00003",X"FFC07",X"FFF8F",X"FFF9F",X"E0007",X"FFFFF",
X"FF000",X"00000",X"0003F",X"FFFFF",X"00FFF",X"FFF00",X"00000",X"03FC0",X"3FFFF",X"FFFE0",X"00007",
X"FFFF0",X"03FF0",X"00000",X"000FF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 421
X"00000",X"003EF",X"C0000",X"00000",X"00000",X"00003",X"FFC07",X"FFFFF",X"FFFBF",X"F0007",X"FFFFF",
X"FF000",X"00000",X"0003F",X"FFFFF",X"00FFF",X"FFF00",X"00000",X"03FC0",X"3FFFF",X"FFFE0",X"00007",
X"FFFF0",X"3FFFF",X"00000",X"000FF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 422
X"00000",X"003FF",X"C0000",X"00000",X"00000",X"00003",X"FFC07",X"FFFFF",X"FFFFF",X"F8007",X"FFFFF",
X"FF000",X"00000",X"0003F",X"FFFFF",X"007FF",X"FFF00",X"00000",X"03FC0",X"3FFFF",X"FFFE0",X"00007",
X"FFFF0",X"1FFFF",X"00000",X"000FF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 423
X"00000",X"003FF",X"C0000",X"00000",X"00000",X"00003",X"FFC07",X"FFFFF",X"FFFFF",X"F8007",X"FFFFF",
X"FF000",X"00000",X"0003F",X"FFFFF",X"007FF",X"FFF1E",X"00000",X"03FDF",X"FFFFF",X"FFFE0",X"00007",
X"FFFF0",X"1FFFF",X"00000",X"01FFF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 424
X"00000",X"003FF",X"E0000",X"00000",X"00000",X"00003",X"FFC07",X"FFFFF",X"FFFFF",X"FD007",X"FFFFF",
X"FF000",X"00000",X"0003F",X"FFFFF",X"007FF",X"FFF1E",X"00000",X"03FDF",X"FFFFF",X"FFFF0",X"00007",
X"FFFF0",X"1FFFF",X"00000",X"01FFF",X"FFFFF",X"FE000",X"00000",X"00000",X"00000",X"00000",-- row 425
X"00000",X"003FF",X"E0000",X"00000",X"00000",X"00003",X"FFC07",X"FFFFF",X"FFFFF",X"FF007",X"FFFFF",
X"FF800",X"00000",X"0003F",X"FFFFF",X"007FF",X"FFF1E",X"00000",X"03FDF",X"FFFFF",X"FFFF0",X"00007",
X"FFFF0",X"1FFFF",X"00000",X"01FFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 426
X"00000",X"001FF",X"E0000",X"00000",X"00000",X"00003",X"FFC07",X"FFFFF",X"FFFFF",X"FF807",X"FFFFF",
X"FF800",X"00000",X"0003F",X"FFFFF",X"007FF",X"FFF3E",X"00000",X"03FDF",X"FFFFF",X"FFFF0",X"C0007",
X"FFFFF",X"FFFFF",X"00000",X"0FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 427
X"00000",X"001FF",X"F8000",X"00000",X"00000",X"00003",X"FFC07",X"FFFFF",X"FFFFF",X"FF807",X"FFFFF",
X"FF800",X"00000",X"0003F",X"FFFFF",X"007FF",X"FFF3F",X"C0000",X"03FDF",X"FFFFF",X"FFFFF",X"FE007",
X"FFFFF",X"FFFFF",X"00000",X"0FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 428
X"00000",X"000FF",X"F8000",X"00000",X"00000",X"00003",X"FFC07",X"FFFFF",X"FFFFF",X"FF807",X"FFFFF",
X"FFC00",X"00000",X"0003F",X"FFFFF",X"007FF",X"FFF3F",X"C07F0",X"03FDF",X"FFFFF",X"FFFFF",X"FE20F",
X"FFFFF",X"FFFFF",X"01F00",X"3FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 429
X"00000",X"000FF",X"FC000",X"00000",X"00000",X"00003",X"FFC07",X"FFFFF",X"FFFFF",X"FF807",X"FFFFF",
X"FFC00",X"00000",X"0003F",X"FFFFF",X"007FF",X"FFF3F",X"C07FF",X"FFFFF",X"FFFFF",X"FFFFF",X"FE20F",
X"FFFFF",X"FFFFF",X"FFF00",X"3FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 430
X"00000",X"000FF",X"FC000",X"00000",X"00000",X"00003",X"FFC07",X"FFFFF",X"FFFFF",X"FF807",X"FFFFF",
X"FFE00",X"00000",X"0003F",X"FFFFF",X"E47FF",X"FFF3F",X"C27FF",X"FFFFF",X"FFFFF",X"FFFFF",X"FE20F",
X"FFFFF",X"FFFFF",X"FFFF0",X"3FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 431
X"00000",X"000FF",X"FC600",X"00000",X"00000",X"00003",X"FFC07",X"FFFFF",X"FFFFF",X"FFC07",X"FFFFF",
X"FFE00",X"00000",X"0003F",X"FFFFF",X"E47FF",X"FFF3F",X"C47FF",X"FFFFF",X"FFFFF",X"FFFFF",X"FE21F",
X"FFFFF",X"FFFFF",X"FFFF0",X"3FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 432
X"00000",X"000FF",X"FF780",X"00000",X"00000",X"00003",X"FFC07",X"FFFFF",X"FFFFF",X"FFC07",X"FFFFF",
X"FFF00",X"00000",X"0003F",X"FFFFF",X"E67FF",X"FFF3F",X"C47FF",X"FFFFF",X"FFFFF",X"FFFFF",X"FE27F",
X"FFFFF",X"FFFFF",X"FFFF0",X"3FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 433
X"00000",X"0007F",X"FFF80",X"00000",X"00000",X"00003",X"FFC0F",X"FFFFF",X"FFFFF",X"FFC07",X"FFFFF",
X"FFF00",X"06C00",X"6003F",X"FFFFF",X"EE7FF",X"FFF3F",X"C4FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF77F",
X"FFFFF",X"FFFFF",X"FFFF0",X"3FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 434
X"00000",X"000FF",X"FFF00",X"00000",X"00000",X"00003",X"FFFFF",X"FFFFF",X"FFFFF",X"FFDE7",X"FFFFF",
X"FFF0F",X"FFF00",X"F803F",X"FFFFF",X"FFFFF",X"FFFBF",X"FCFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFF0",X"3FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 435
X"00000",X"000FF",X"FFF80",X"00000",X"3FFF8",X"00003",X"FFFFF",X"FFFFF",X"FFFFF",X"FFDFF",X"FFFFF",
X"FFF0F",X"FFF0C",X"F803F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFF0",X"3FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 436
X"00000",X"001FF",X"FFF00",X"00000",X"3FFF8",X"00003",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFF0F",X"FFF0D",X"FC03F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFF0",X"3FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 437
X"00000",X"001FF",X"FFF00",X"00000",X"3FFF8",X"00003",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFF0F",X"FFF0F",X"FE03F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFF0",X"3FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 438
X"00000",X"001FF",X"FFE00",X"00000",X"3FFF8",X"00043",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFF0F",X"FFF7F",X"FE03F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFF0",X"3FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 439
X"00000",X"001FF",X"FFC00",X"00000",X"7FFFC",X"00043",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFF0F",X"FFF7F",X"FF03F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFF0",X"3FFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 440
X"00000",X"000FF",X"FFC00",X"00000",X"7FFFE",X"00043",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFF0F",X"FFF7F",X"FF83F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 441
X"00000",X"000FF",X"FFC00",X"00030",X"7FFFE",X"000C3",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFF0F",X"FFF7F",X"FF83F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 442
X"00000",X"000FF",X"FFC00",X"0003E",X"7FFFE",X"000E3",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFF0F",X"FFF7F",X"FF83F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 443
X"00000",X"000FF",X"FF800",X"00E3E",X"7FFFE",X"600EF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFF0F",X"FFF7F",X"FF81F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF000",X"00000",X"00000",X"00000",X"00000",-- row 444
X"00000",X"000FF",X"FF000",X"00FFE",X"7FFFE",X"798EF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFF0F",X"FFF7F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF000",X"00008",X"00000",X"00000",X"00000",-- row 445
X"00000",X"000FF",X"FE000",X"00FFE",X"7FFFE",X"798EF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFF0F",X"FFF7F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF000",X"006FC",X"00000",X"00000",X"00000",-- row 446
X"00000",X"000FF",X"FF000",X"00FFF",X"FFFFE",X"F98EF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFF0F",X"FFF7F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF000",X"5FFFE",X"00000",X"00000",X"00000",-- row 447
X"00000",X"000FF",X"FF000",X"00FFF",X"FFFFF",X"FFFEF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFCF",X"FFF7F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF005",X"0FFFD",X"00000",X"00000",X"00000",-- row 448
X"00000",X"000FF",X"FF000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFCF",X"FFF7F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF050",X"07FFD",X"00000",X"00000",X"00000",-- row 449
X"00000",X"000FF",X"FF000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFCF",X"FFF7F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF500",X"2FFFC",X"80000",X"00000",X"00000",-- row 450
X"00000",X"0007F",X"FF000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFCF",X"FFF7F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF002",X"87FFC",X"80000",X"00000",X"00000",-- row 451
X"00000",X"0007F",X"FF000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFCF",X"FFF7F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF028",X"07FBC",X"40000",X"00000",X"00000",-- row 452
X"00000",X"000FF",X"FF000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFDF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFA80",X"0739C",X"20000",X"00000",X"00000",-- row 453
X"00000",X"000FF",X"FF000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFDF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF000",X"0739C",X"00000",X"00000",X"00000",-- row 454
X"00000",X"0007F",X"FF000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF000",X"073DC",X"10000",X"00000",X"00000",-- row 455
X"00000",X"000FF",X"FF000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFE00",X"073BC",X"08000",X"00000",X"00000",-- row 456
X"00000",X"000FF",X"FE000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFC0",X"0739C",X"04000",X"00000",X"00000",-- row 457
X"00000",X"000FF",X"FE000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFF8",X"0739C",X"00000",X"00000",X"00000",-- row 458
X"00000",X"000FF",X"FE000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"0739E",X"02000",X"00000",X"00000",-- row 459
X"00000",X"000FF",X"FE000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"E739D",X"01000",X"00000",X"00000",-- row 460
X"00000",X"000FF",X"FE000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF79C",X"80800",X"00000",X"00000",-- row 461
X"00000",X"0007F",X"FE000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFDE",X"40400",X"00000",X"00000",-- row 462
X"00000",X"0007F",X"FE000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF01F",X"FFFFE",X"10200",X"00000",X"00000",-- row 463
X"00000",X"000FF",X"FE000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF000",X"1FFFF",X"FC19E",X"00000",X"00000",-- row 464
X"00000",X"0007F",X"FE000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF000",X"0FFFF",X"FFC54",X"00000",X"00000",-- row 465
X"00000",X"0007F",X"FE000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF000",X"0FFFE",X"03FBC",X"00000",X"00000",-- row 466
X"00000",X"0007F",X"FE000",X"00FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF004",X"0FFFE",X"001F4",X"00000",X"00000",-- row 467
X"00000",X"001FF",X"FE000",X"03FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FF004",X"FFFFE",X"0003E",X"00000",X"00000",-- row 468
X"00000",X"00FFF",X"FF000",X"07FFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFE",X"0011F",X"00000",X"00000",-- row 469
X"00000",X"00FFF",X"FF000",X"1FFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFBFF",X"FFF80",X"00000",-- row 470
X"00000",X"00FFF",X"FF807",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFF8",X"00000",-- row 471
X"00000",X"01FFF",X"FF81F",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFE",X"00000",-- row 472
X"00000",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFE",X"00000",X"00000",X"00000",-- row 473
X"00000",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFE",X"00000",X"00000",X"00000",-- row 474
X"00000",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFE",X"00000",X"00000",X"00000",-- row 475
X"00000",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"E0000",X"00000",X"00000",-- row 476
X"00000",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FC000",X"00000",X"00000",-- row 477
X"00000",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFC00",X"00000",X"00000",-- row 478
X"00000",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",
X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFFFF",X"FFF00",X"00000",X"00000",-- row 479
others=>X"00000");

begin

address <= unsigned(row(8 downto 0)) & word_col;
ncol <= to_integer(unsigned(next_col));

process(clk)
begin 
	if rising_edge(clk) then
		mem_out <= unsigned(framebuffer(to_integer(address))); --fill with zeros?
	end if;
end process;


process(ncol)
begin
	word_col <= "00000";
	load <= false;
	if ncol = 831 then
		word_col <= "00000";
	elsif ncol = 0 then
		load <= true;
	else 
		for i in 1 to 31 loop
			if ncol = i *20 -1 then 
				word_col <= to_unsigned(i, word_col'length);
			elsif ncol = i * 20 then
				load <= true;
			end if;
		end loop;
	end if;
end process;



process(clk) --shift register
begin
	if rising_edge(clk) then
		if load then
			pixel_vec <= mem_out;
		else 
			pixel_vec <= pixel_vec(18 downto 0) & '0';
		end if;
	end if;
end process;

pixel <= pixel_vec(19);
			
			


end Behavioral;

